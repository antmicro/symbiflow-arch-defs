module top(
    input wire in,
    output wire out
);

(* keep, LOC="GTPE2_CHANNEL_X0Y0" *)
GTPE2_CHANNEL #(
            .ACJTAG_RESET(1'b0),
            .ACJTAG_DEBUG_MODE(1'b0),
            .ACJTAG_MODE(1'b0),
            .UCODEER_CLR(1'b0),
            .RXBUFRESET_TIME(5'b01100),
            .RXCDRPHRESET_TIME(5'b10110),
            .RXCDRFREQRESET_TIME(5'b10011),
            .RXPMARESET_TIME(5'b10001),
            .RXPCSRESET_TIME(5'b11010),
            .RXLPMRESET_TIME(7'b0010100),
            .RXISCANRESET_TIME(5'b10111),
            .RXSYNC_OVRD(1'b1),
            .TXSYNC_OVRD(1'b1),
            .RXSYNC_SKIP_DA(1'b0),
            .TXSYNC_SKIP_DA(1'b1),
            .TXSYNC_MULTILANE(1'b0),
            .RXSYNC_MULTILANE(1'b0),
            .TXPCSRESET_TIME(5'b10001),
            .TXPMARESET_TIME(5'b01111),
            .RX_XCLK_SEL("RXUSR"),
            .RX_DATA_WIDTH(40),
            .RX_CLK25_DIV(15),
            .RX_CM_SEL(2'b01),
            .RXPRBS_ERR_LOOPBACK(1'b1),
            .SATA_BURST_SEQ_LEN(4'b0001),
            .OUTREFCLK_SEL_INV(2'b11),
            .SATA_BURST_VAL(3'b000),
            .RXOOB_CFG(7'b1011001),
            .SAS_MIN_COM(49),
            .SATA_MIN_BURST(17),
            .SATA_EIDLE_VAL(3'b110),
            .SATA_MIN_WAKE(15),
            .SATA_MIN_INIT(58),
            .SAS_MAX_COM(86),
            .SATA_MAX_BURST(44),
            .SATA_MAX_WAKE(5),
            .SATA_MAX_INIT(30),
            .RXOSCALRESET_TIMEOUT(5'b00110),
            .RXOSCALRESET_TIME(5'b00111),
            .TRANS_TIME_RATE(8'b11001010),
            .PMA_LOOPBACK_CFG(1'b1),
            .TX_PREDRIVER_MODE(1'b0),
            .TX_EIDLE_DEASSERT_DELAY(3'b010),
            .TX_EIDLE_ASSERT_DELAY(3'b111),
            .TX_LOOPBACK_DRIVE_HIZ("TRUE"),
            .TX_DRIVE_MODE("DIRECT"),
            .PD_TRANS_TIME_TO_P2(8'b01010011),
            .PD_TRANS_TIME_NONE_P2(8'b01000110),
            .PD_TRANS_TIME_FROM_P2(12'b011100101011),
            .PCS_PCIE_EN("TRUE"),
            .TXBUF_RESET_ON_RATE_CHANGE("TRUE"),
            .TXBUF_EN("FALSE"),
            .TXGEARBOX_EN("FALSE"),
            .GEARBOX_MODE(3'b011),
            .RXLPM_HOLD_DURING_EIDLE(1'b1),
            .RX_OS_CFG(13'b1010101001000),
            .RXLPM_LF_CFG(18'b110000110011111000),
            .RXLPM_HF_CFG(14'b01111001010101),
            .ES_QUALIFIER(80'b10111110101011001100110001000100110110010011011010100001011101100001100000001110),
            .ES_QUAL_MASK(80'b00111111111101101101001110000110110101101011001011110101110010010111011010111000),
            .ES_SDATA_MASK(80'b01101011000011111101111101100110110010001110101110110010111001110011001100010001),
            .ES_PRESCALE(5'b00001),
            .ES_VERT_OFFSET(9'b000011100),
            .ES_HORZ_OFFSET(12'b101101011100),
            .RX_DISPERR_SEQ_MATCH("FALSE"),
            .DEC_PCOMMA_DETECT("TRUE"),
            .DEC_MCOMMA_DETECT("TRUE"),
            .DEC_VALID_COMMA_ONLY("TRUE"),
            .ES_ERRDET_EN("TRUE"),
            .ES_EYE_SCAN_EN("FALSE"),
            .ES_CONTROL(6'b001011),
            .ALIGN_COMMA_ENABLE(10'b0011110000),
            .ALIGN_MCOMMA_VALUE(10'b1110110001),
            .RXSLIDE_MODE("PCS"),
            .ALIGN_PCOMMA_VALUE(10'b0010000011),
            .ALIGN_COMMA_WORD(2),
            .RX_SIG_VALID_DLY(23),
            .ALIGN_PCOMMA_DET("FALSE"),
            .ALIGN_MCOMMA_DET("FALSE"),
            .SHOW_REALIGN_COMMA("TRUE"),
            .ALIGN_COMMA_DOUBLE("TRUE"),
            .RXSLIDE_AUTO_WAIT(6),
            .CLK_CORRECT_USE("FALSE"),
            .CLK_COR_SEQ_1_ENABLE(4'b0011),
            .CLK_COR_SEQ_1_1(10'b0001110010),
            .CLK_COR_MAX_LAT(8),
            .CLK_COR_SEQ_1_2(10'b1000111110),
            .CLK_COR_MIN_LAT(27),
            .CLK_COR_SEQ_1_3(10'b1101001001),
            .CLK_COR_REPEAT_WAIT(28),
            .CLK_COR_SEQ_1_4(10'b0101100011),
            .CLK_COR_SEQ_2_USE("TRUE"),
            .CLK_COR_SEQ_2_ENABLE(4'b1011),
            .CLK_COR_SEQ_2_1(10'b1000111010),
            .CLK_COR_KEEP_IDLE("TRUE"),
            .CLK_COR_PRECEDENCE("FALSE"),
            .CLK_COR_SEQ_LEN(4),
            .CLK_COR_SEQ_2_2(10'b0111111100),
            .CLK_COR_SEQ_2_3(10'b1011000011),
            .RXGEARBOX_EN("FALSE"),
            .CLK_COR_SEQ_2_4(10'b0110110111),
            .CHAN_BOND_SEQ_1_ENABLE(4'b0101),
            .CHAN_BOND_SEQ_1_1(10'b0100101011),
            .CHAN_BOND_SEQ_LEN(1),
            .CHAN_BOND_SEQ_1_2(10'b1010110001),
            .CHAN_BOND_KEEP_ALIGN("TRUE"),
            .CHAN_BOND_SEQ_1_3(10'b0011100111),
            .CHAN_BOND_SEQ_1_4(10'b1111010100),
            .CHAN_BOND_SEQ_2_ENABLE(4'b1000),
            .CHAN_BOND_SEQ_2_USE("TRUE"),
            .CHAN_BOND_SEQ_2_1(10'b0010101001),
            .FTS_LANE_DESKEW_CFG(4'b1101),
            .FTS_LANE_DESKEW_EN("FALSE"),
            .CHAN_BOND_SEQ_2_2(10'b0001001000),
            .FTS_DESKEW_SEQ_ENABLE(4'b0100),
            .CBCC_DATA_SOURCE_SEL("DECODED"),
            .CHAN_BOND_SEQ_2_3(10'b0100100000),
            .CHAN_BOND_MAX_SKEW(10),
            .CHAN_BOND_SEQ_2_4(10'b0110000001),
            .RXDLY_TAP_CFG(16'b1010001110010010),
            .RXDLY_CFG(16'b0100011111000101),
            .RXPH_MONITOR_SEL(5'b10001),
            .RX_DDI_SEL(6'b110011),
            .TX_XCLK_SEL("TXOUT"),
            .RXBUF_EN("FALSE"),
            .TXOOB_CFG(1'b0),
            .LOOPBACK_CFG(1'b0),
            .TXPI_CFG5(3'b000),
            .TXPI_CFG4(1'b1),
            .TXPI_CFG3(1'b0),
            .TXPI_CFG2(2'b11),
            .TXPI_CFG1(2'b11),
            .TXPI_CFG0(2'b01),
            .SATA_PLL_CFG("VCO_1500MHZ"),
            .TXPHDLY_CFG(24'b011001100011111101011100),
            .TXDLY_CFG(16'b0001001111000001),
            .TXDLY_TAP_CFG(16'b0100110011010010),
            .TXPH_CFG(16'b0100011100111001),
            .TXPH_MONITOR_SEL(5'b00000),
            .RX_BIAS_CFG(16'b1001111011010001),
            .RXOOB_CLK_CFG("FABRIC"),
            .TX_CLKMUX_EN(1'b1),
            .RX_CLKMUX_EN(1'b0),
            .TERM_RCAL_CFG(15'b011011000110000),
            .TERM_RCAL_OVRD(3'b101),
            .TX_CLK25_DIV(12),
            .PMA_RSV5(1'b0),
            .PMA_RSV4(4'b0010),
            .TX_DATA_WIDTH(20),
            .PCS_RSVD_ATTR(48'b101010101110110011011101010011001001001100110010),
            .TX_MARGIN_FULL_1(7'b0000001),
            .TX_MARGIN_FULL_0(7'b0110001),
            .TX_MARGIN_FULL_3(7'b1000011),
            .TX_MARGIN_FULL_2(7'b1100011),
            .TX_MARGIN_LOW_0(7'b0001101),
            .TX_MARGIN_FULL_4(7'b1100110),
            .TX_MARGIN_LOW_2(7'b1001000),
            .TX_MARGIN_LOW_1(7'b1010111),
            .TX_MARGIN_LOW_4(7'b0010000),
            .TX_MARGIN_LOW_3(7'b0001000),
            .TX_DEEMPH1(6'b110001),
            .TX_DEEMPH0(6'b011000),
            .TX_RXDETECT_REF(3'b000),
            .TX_MAINCURSOR_SEL(1'b1),
            .PMA_RSV3(2'b00),
            .PMA_RSV7(1'b1),
            .PMA_RSV6(1'b0),
            .TX_RXDETECT_CFG(14'b11010010110011),
            .CLK_COMMON_SWING(1'b1),
            .RX_CM_TRIM(4'b0110),
            .RXLPM_CFG1(1'b1),
            .RXLPM_CFG(4'b1110),
            .PMA_RSV2(32'b10110101001111001100010110000111),
            .DMONITOR_CFG(24'b100001101001000011010010),
            .RXLPM_BIAS_STARTUP_DISABLE(1'b1),
            .RXLPM_HF_CFG3(4'b0100),
            .TXOUT_DIV(4),
            .RXOUT_DIV(8),
            .CFOK_CFG(43'b0000110001101010101100111110110010011000010),
            .CFOK_CFG3(7'b0110110),
            .RXPI_CFG0(3'b100),
            .RXLPM_CM_CFG(1'b0),
            .CFOK_CFG5(2'b11),
            .RXLPM_LF_CFG2(5'b00011),
            .RXLPM_HF_CFG2(5'b10101),
            .RXLPM_IPCM_CFG(1'b0),
            .RXLPM_INCM_CFG(1'b0),
            .CFOK_CFG4(1'b0),
            .CFOK_CFG6(4'b1000),
            .RXLPM_GC_CFG(9'b001110100),
            .RXLPM_GC_CFG2(3'b110),
            .RXPI_CFG1(1'b0),
            .RXPI_CFG2(1'b1),
            .RXLPM_OSINT_CFG(3'b101),
            .ES_CLK_PHASE_SEL(1'b0),
            .USE_PCS_CLK_PHASE_SEL(1'b1),
            .CFOK_CFG2(7'b1000111),
            .ADAPT_CFG0(20'b10111011010101001111),
            .TXPI_PPM_CFG(8'b11001001),
            .TXPI_GREY_SEL(1'b1),
            .TXPI_INVSTROBE_SEL(1'b1),
            .TXPI_PPMCLK_SEL("TXUSRCLK"),
            .TXPI_SYNFREQ_PPM(3'b101),
            .TST_RSV(32'b00101001001011100000001000110101),
            .PMA_RSV(32'b00101010100101011101011000011011),
            .RX_BUFFER_CFG(6'b000001),
            .RXBUF_THRESH_OVRD("FALSE"),
            .RXBUF_RESET_ON_EIDLE("TRUE"),
            .RXBUF_THRESH_UNDFLW(44),
            .RXBUF_EIDLE_HI_CNT(4'b1011),
            .RXBUF_EIDLE_LO_CNT(4'b0011),
            .RXBUF_ADDR_MODE("FAST"),
            .RXBUF_THRESH_OVFLW(1),
            .RX_DEFER_RESET_BUF_EN("TRUE"),
            .RXBUF_RESET_ON_COMMAALIGN("TRUE"),
            .RXBUF_RESET_ON_RATE_CHANGE("TRUE"),
            .RXBUF_RESET_ON_CB_CHANGE("TRUE"),
            .TXDLY_LCFG(9'b100001011),
            .RXDLY_LCFG(9'b100101011),
            .RXPH_CFG(24'b111011000011011001001110),
            .RXPHDLY_CFG(24'b011100111010101011111001),
            .RX_DEBUG_CFG(14'b11100111111000),
            .ES_PMA_CFG(10'b1000110010),
            .RXCDR_PH_RESET_ON_EIDLE(1'b1),
            .RXCDR_FR_RESET_ON_EIDLE(1'b0),
            .RXCDR_HOLD_DURING_EIDLE(1'b1),
            .RXCDR_LOCK_CFG(6'b010011),
            .RXCDR_CFG(83'b11011011100001110001001101000010110010000001101010000011010111001011010011100111111),
            .IS_TXUSRCLK_INVERTED(1),
            .IS_TXUSRCLK2_INVERTED(0),
            .IS_TXPHDLYTSTCLK_INVERTED(1),
            .IS_SIGVALIDCLK_INVERTED(1),
            .IS_RXUSRCLK_INVERTED(0),
            .IS_RXUSRCLK2_INVERTED(0),
            .IS_DRPCLK_INVERTED(1),
            .IS_DMONITORCLK_INVERTED(0),
            .IS_CLKRSVD0_INVERTED(0),
            .IS_CLKRSVD1_INVERTED(0)
    ) gtp_channel_0 (
            .DRPCLK(in),
	    .DRPRDY(out)
    );
endmodule
