(* whitebox *)
(* MODEL_NAME="GND" *)
module GND_CELL (
    output wire GND
);

    assign GND = 1'b0;

endmodule
