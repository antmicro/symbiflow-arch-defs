(* whitebox *)
module DELAY (
	IN,
	OUT
);

input wire IN;
output wire OUT;

assign OUT = IN;

endmodule
