module top(
    input wire in,
    output wire out
);

(* keep, LOC="GTPE2_COMMON_X0Y0" *)
GTPE2_COMMON #(
            .PLL0_CFG(27'b001011100100001101100001010),
            .PLL0_REFCLK_DIV(1),
            .PLL0_FBDIV_45(5),
            .PLL0_FBDIV(1),
            .PLL0_LOCK_CFG(9'b100010110),
            .PLL0_INIT_CFG(24'b110100010100101001101100),
            .RSVD_ATTR0(16'b0100101010100101),
            .PLL1_DMON_CFG(1'b0),
            .PLL0_DMON_CFG(1'b0),
            .COMMON_CFG(32'b10010001111100110111001011011010),
            .PLL_CLKOUT_CFG(8'b11011111),
            .BIAS_CFG(64'b0000110100110111011100001111100100110010001111100001111111111111),
            .RSVD_ATTR1(16'b0010110110111111),
            .PLL1_INIT_CFG(24'b100001100010100010111101),
            .PLL1_LOCK_CFG(9'b001110000),
            .PLL1_REFCLK_DIV(1),
            .PLL1_FBDIV_45(4),
            .PLL1_FBDIV(3),
            .PLL1_CFG(27'b111010010111111101110000010),
            .IS_GTGREFCLK1_INVERTED(0),
            .IS_GTGREFCLK0_INVERTED(1),
            .IS_PLL0LOCKDETCLK_INVERTED(1),
            .IS_PLL1LOCKDETCLK_INVERTED(1),
            .IS_DRPCLK_INVERTED(1)
) GTPE2_COMMON_X0Y0 (
        .GTREFCLK0(in),
	.PLL0OUTCLK(out)
    );
endmodule
