(* whitebox *)
(* MODEL_NAME="VCC" *)
module VCC_CELL (
    output wire VCC
);

    assign VCC = 1'b1;

endmodule
